
module pkt_ctrler #() (
    // General I/O
    input   logic                                       clk,
    input   logic                                       rst,

    input   logic                                       in_enque_en,
    output  logic                                       in_valid,
    
    input   logic                                       out_deque_en,
    output  logic                                       out_valid,
);


endmodule